library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_unsigned.all;



entity pipeline is
port(
    reset, clock : in std_logic --pinos do reset e do clock para o PC
);
end entity;


architecture behavior of pipeline is

      -- PC e MUXES para o PC
     signal PC : std_logic_vector (7 downto 0); --sinal para o PC
     signal pc_next : std_logic_vector(7 downto 0);
     signal pc_branch_end : std_logic_vector(7 downto 0);
     signal branch_taken : std_logic; -- sinal para indicar se o branch e tomado ou nao


     signal decode_opcode : std_logic_vector(3 downto 0);

     -- MEMORIA DE INSTRU�AO
     type memoria_inst_t is array (integer range 0 to 255) of std_logic_vector (19 downto 0);
     signal memoria_instrucoes       : memoria_inst_t;
     signal memoria_instrucoes_out   : std_logic_vector (19 downto 0);



    -- MEMORIA DE DADOS (cada posi��o 16 bits)
    type memoria_dados_t is array (integer range 0 to 255) of std_logic_vector (15 downto 0);
    signal memoria_dados       : memoria_dados_t;
    signal memoria_dados_out   : std_logic_vector (15 downto 0); -- valor
    signal endereco_mem        : std_logic_vector (15 downto 0);

    -- BANCO DE REGISTRADORES DO MIPS
    type registradores is array (integer range 0 to 15) of std_logic_vector(15 downto 0); -- indices sendo representador por inteiros por isso a conversao
    signal banco_reg : registradores;

  


     -- EST�GIO IF/ID
    signal IF_ID_PC : std_logic_vector(7 downto 0);
    signal IF_ID_instruction : std_logic_vector(19 downto 0);
    
    -- EST�GIO ID/EX
    signal ID_EX_opcode : std_logic_vector(3 downto 0);
    signal ID_EX_reg_rs, ID_EX_reg_rt, ID_EX_reg_rd : std_logic_vector(3 downto 0);
    signal ID_EX_valor_rs, ID_EX_valor_rt : std_logic_vector(15 downto 0);
    signal ID_EX_imediato : std_logic_vector(7 downto 0);
    
    -- EST�GIO EX/MEM
    signal EX_MEM_opcode : std_logic_vector(3 downto 0);
    signal EX_MEM_resultado_ula : std_logic_vector(15 downto 0);
    signal EX_MEM_valor_rt : std_logic_vector(15 downto 0);
    signal EX_MEM_reg_dest : std_logic_vector(3 downto 0);
    
    -- EST�GIO MEM/WB
    signal MEM_WB_opcode : std_logic_vector(3 downto 0);
    signal MEM_WB_resultado_ula : std_logic_vector(15 downto 0);
    signal MEM_WB_dado_mem : std_logic_vector(15 downto 0);
    signal MEM_WB_reg_dest : std_logic_vector(3 downto 0);

   

begin

    -- buscar instru��o
    memoria_instrucoes_out <= memoria_instrucoes(conv_integer(PC)) when reset = '0' else
    (others => '0');

    -- buscar dados da memoria
    memoria_dados_out <= memoria_dados(conv_integer(endereco_mem(7 downto 0)));
  
    -- logica para o PC	
    pc_next <= pc_branch_end when branch_taken = '1' else
               PC + 1;



  

    process(reset, clock)
    begin
        if reset = '1' then
            PC <= (others => '0');
            banco_reg <= (others => (others => '0')); -- limpa todos no reset
            memoria_dados <= (others => (others => '0'));  -- limpa mem�ria de dados
	    memoria_instrucoes <= (others => (others => '0'));
	    IF_ID_PC <= (others => '0');
	    IF_ID_instruction <= (others => '0');
	    ID_EX_opcode <= (others => '0');

	    		-------------------***/ INSTRU�OES \***-------------------


	              -- TIPO I: | OPCODE(4) | RT(4) | RS(4) | IMD(8)| banco_reg(rt) <- imd    
	memoria_instrucoes(0) <= "01000010000000001010"; -- LDI banco_reg(2) <- 10
        memoria_instrucoes(1) <= "01000011000000001010"; -- LDI banco_reg(3) <- 10
	memoria_instrucoes(2) <= "01001010000000000101"; -- LDI banco_reg(10)<- 5
	memoria_instrucoes(3) <= "01001011000000000010"; -- LDI banco_reg(11)<- 2
		      
		      -- TIPO R: | OPCODE(4) | RD(4) | RS(4) | RT(4) | don't care(4)| banco_reg(rd) <- rs + rt
	memoria_instrucoes(4) <= "00010100001000110000"; -- ADD banco_reg(4) <-banco_reg(2) + banco_reg(3) |10 + 10| 
        memoria_instrucoes(5) <= "00100101001010100000"; -- SUB banco_reg(5) <- banco_reg(2) - banco_reg(10) | 10 - 5|
        memoria_instrucoes(6) <= "00110110101110100000"; -- MUL banco_reg(6) <- banco_reg(11) * banco_reg(10) | 2 * 5|     

	               -- TIPO I: | OPCODE(4) | RT(4) | RS(4) | IMD(8)| banco_reg(rt) <- banco_reg(rs) + imd
	memoria_instrucoes(7) <= "01010111101100000010"; -- ADDI banco_reg(7) <- banco_reg(11) + 2  | 2 + 2 |		
 	memoria_instrucoes(8) <= "01101000001100001001"; -- SUBI banco_reg(8) <- banco_reg(3) - 9 | 10 - 9 |
	memoria_instrucoes(9) <= "01111001101100000100"; -- MULI banco_reg(9) <- banco_reg(11) * 5 | 2 * 5| -- ANALISAR DEPOIS
			-- SW Mem[rs + imd] <- rt
	memoria_instrucoes(10) <= "10011000000000000100"; -- SW mem_dados(4) <- banco_reg(rt-8)|1| 
	memoria_instrucoes(12) <= "10010010000000001010";  -- SW mem_dados(10) <- banco_reg(rt-2)|10|
			-- LW rt <- Mem[rs + imd]
	memoria_instrucoes(13) <= "10001100000000000100"; -- LW banco_reg(12) <- mem_dados(4)|1|
	memoria_instrucoes(14) <= "10001101000000001010"; -- LW banco_reg(13) <- mem_dados(10)|10|
			-- Formato J: JMP ( OPCODE(4) | ENDERECO(8) | 00000000)
	memoria_instrucoes(15) <= "10100011001000000000"; -- PC <- END 50

		        --Formato B:  (OPCODE(4) | RS(4) | RT(4) | DESLOC(8)
	memoria_instrucoes(50) <= "10111101101000110010"; -- BEQ reg(12)|10| == reg(10)|5| pc<= 100
	memoria_instrucoes(51) <= "00101101110111000000"; -- SUB reg(12) <- 10 - 1 
	memoria_instrucoes(52) <= "10100011001000000000"; -- PC <- END 50
	
	

			-------------------***/ INSTRU�OES \***-------------------


   elsif  clock'event and clock = '1' then
           
            -- garante r0 = 0 (sempre)
            banco_reg(0) <= (others => '0');


	    --------------------------------
            -- EST�GIO IF (Instruction Fetch)
            --------------------------------
	    PC <= pc_next;


	    ------------- IF -> ID -------------
	    IF_ID_PC <= PC; -- recebe PC
	    IF_ID_instruction <= memoria_instrucoes_out;  --IF recebe memoria de instrucao



	    --------------------------------
            -- EST�GIO ID (Instruction Decode)
            --------------------------------
	    decode_opcode <= IF_ID_instruction(19 downto 16);
	
	    -- ID -> EX
	    ID_EX_opcode <= decode_opcode;
	    ID_EX_reg_rs <= IF_ID_instruction(15 downto 12);
	    ID_EX_reg_rt <= IF_ID_instruction(11 downto 8);
	    ID_EX_reg_rd <= IF_ID_instruction(7 downto 4);
	    ID_EX_imediato <= IF_ID_instruction(7 downto 0);
	    
	    ID_EX_valor_rs <= banco_reg(conv_integer(ID_EX_reg_rs));
	    ID_EX_valor_rt <= banco_reg(conv_integer(ID_EX_reg_rt));


	    --------------------------------
            -- EST�GIO EX (Execute)
            --------------------------------
		

	     --ADD	
	    if ID_EX_opcode = "0001" then
	     EX_MEM_resultado_ula <= ID_EX_valor_rs + ID_EX_valor_rt;
	    end if;


	    -- EX -> MEM
	    EX_MEM_opcode <= ID_EX_opcode;
	    EX_MEM_reg_dest <= ID_EX_reg_rd;
		

	    --------------------------------
            -- EST�GIO MEM (Memory Access)
            --------------------------------

	    if EX_MEM_opcode = "1000" then
	    
		MEM_WB_dado_mem <= memoria_dados(conv_integer(EX_MEM_resultado_ula(7 downto 0)));
	    end if;

	
	
	    -- MEM -> WB
	    MEM_WB_opcode <= EX_MEM_opcode;
	    MEM_WB_resultado_ula <= EX_MEM_resultado_ula;
	    MEM_WB_reg_dest <= EX_MEM_reg_dest;



	    --------------------------------
            -- EST�GIO WB (Write Back)
            --------------------------------

	    if MEM_WB_opcode = "0001" then  -- ADD
	       if MEM_WB_reg_dest /= "0000" then
	        banco_reg(conv_integer(MEM_WB_reg_dest)) <= MEM_WB_resultado_ula;
	       end if;
	    end if;
	


           end if;
    end process;




end architecture;

